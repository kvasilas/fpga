-- D flip flop rising edge
-- VHDL code
-- https://www.fpga4student.com/2017/02/vhdl-code-for-d-flip-flop.html
library IEEE;
USE IEEE.Std_logic_1164.all;
